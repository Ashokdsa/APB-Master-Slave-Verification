parameter N = 2;
