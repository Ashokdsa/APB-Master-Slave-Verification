`include "seq_item.sv"
